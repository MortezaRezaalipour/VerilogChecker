module top(a, b, c);
input [4:0]a;
input [4:0]b;
output [9:0]c;
assign c = a * b;
endmodule
