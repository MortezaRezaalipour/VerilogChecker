module abs_diff_i8_o4_tb;
reg [7:0] pi;
wire [3:0] po;
abs_diff_i8_o4 dut (pi[7], pi[6], pi[5], pi[4], pi[3], pi[2], pi[1], pi[0], po[3], po[2], po[1], po[0]);
initial
begin
#1 pi=8'b00000000;
#1 $display("%b", po);
#1 pi=8'b00000001;
#1 $display("%b", po);
#1 pi=8'b00000010;
#1 $display("%b", po);
#1 pi=8'b00000011;
#1 $display("%b", po);
#1 pi=8'b00000100;
#1 $display("%b", po);
#1 pi=8'b00000101;
#1 $display("%b", po);
#1 pi=8'b00000110;
#1 $display("%b", po);
#1 pi=8'b00000111;
#1 $display("%b", po);
#1 pi=8'b00001000;
#1 $display("%b", po);
#1 pi=8'b00001001;
#1 $display("%b", po);
#1 pi=8'b00001010;
#1 $display("%b", po);
#1 pi=8'b00001011;
#1 $display("%b", po);
#1 pi=8'b00001100;
#1 $display("%b", po);
#1 pi=8'b00001101;
#1 $display("%b", po);
#1 pi=8'b00001110;
#1 $display("%b", po);
#1 pi=8'b00001111;
#1 $display("%b", po);
#1 pi=8'b00010000;
#1 $display("%b", po);
#1 pi=8'b00010001;
#1 $display("%b", po);
#1 pi=8'b00010010;
#1 $display("%b", po);
#1 pi=8'b00010011;
#1 $display("%b", po);
#1 pi=8'b00010100;
#1 $display("%b", po);
#1 pi=8'b00010101;
#1 $display("%b", po);
#1 pi=8'b00010110;
#1 $display("%b", po);
#1 pi=8'b00010111;
#1 $display("%b", po);
#1 pi=8'b00011000;
#1 $display("%b", po);
#1 pi=8'b00011001;
#1 $display("%b", po);
#1 pi=8'b00011010;
#1 $display("%b", po);
#1 pi=8'b00011011;
#1 $display("%b", po);
#1 pi=8'b00011100;
#1 $display("%b", po);
#1 pi=8'b00011101;
#1 $display("%b", po);
#1 pi=8'b00011110;
#1 $display("%b", po);
#1 pi=8'b00011111;
#1 $display("%b", po);
#1 pi=8'b00100000;
#1 $display("%b", po);
#1 pi=8'b00100001;
#1 $display("%b", po);
#1 pi=8'b00100010;
#1 $display("%b", po);
#1 pi=8'b00100011;
#1 $display("%b", po);
#1 pi=8'b00100100;
#1 $display("%b", po);
#1 pi=8'b00100101;
#1 $display("%b", po);
#1 pi=8'b00100110;
#1 $display("%b", po);
#1 pi=8'b00100111;
#1 $display("%b", po);
#1 pi=8'b00101000;
#1 $display("%b", po);
#1 pi=8'b00101001;
#1 $display("%b", po);
#1 pi=8'b00101010;
#1 $display("%b", po);
#1 pi=8'b00101011;
#1 $display("%b", po);
#1 pi=8'b00101100;
#1 $display("%b", po);
#1 pi=8'b00101101;
#1 $display("%b", po);
#1 pi=8'b00101110;
#1 $display("%b", po);
#1 pi=8'b00101111;
#1 $display("%b", po);
#1 pi=8'b00110000;
#1 $display("%b", po);
#1 pi=8'b00110001;
#1 $display("%b", po);
#1 pi=8'b00110010;
#1 $display("%b", po);
#1 pi=8'b00110011;
#1 $display("%b", po);
#1 pi=8'b00110100;
#1 $display("%b", po);
#1 pi=8'b00110101;
#1 $display("%b", po);
#1 pi=8'b00110110;
#1 $display("%b", po);
#1 pi=8'b00110111;
#1 $display("%b", po);
#1 pi=8'b00111000;
#1 $display("%b", po);
#1 pi=8'b00111001;
#1 $display("%b", po);
#1 pi=8'b00111010;
#1 $display("%b", po);
#1 pi=8'b00111011;
#1 $display("%b", po);
#1 pi=8'b00111100;
#1 $display("%b", po);
#1 pi=8'b00111101;
#1 $display("%b", po);
#1 pi=8'b00111110;
#1 $display("%b", po);
#1 pi=8'b00111111;
#1 $display("%b", po);
#1 pi=8'b01000000;
#1 $display("%b", po);
#1 pi=8'b01000001;
#1 $display("%b", po);
#1 pi=8'b01000010;
#1 $display("%b", po);
#1 pi=8'b01000011;
#1 $display("%b", po);
#1 pi=8'b01000100;
#1 $display("%b", po);
#1 pi=8'b01000101;
#1 $display("%b", po);
#1 pi=8'b01000110;
#1 $display("%b", po);
#1 pi=8'b01000111;
#1 $display("%b", po);
#1 pi=8'b01001000;
#1 $display("%b", po);
#1 pi=8'b01001001;
#1 $display("%b", po);
#1 pi=8'b01001010;
#1 $display("%b", po);
#1 pi=8'b01001011;
#1 $display("%b", po);
#1 pi=8'b01001100;
#1 $display("%b", po);
#1 pi=8'b01001101;
#1 $display("%b", po);
#1 pi=8'b01001110;
#1 $display("%b", po);
#1 pi=8'b01001111;
#1 $display("%b", po);
#1 pi=8'b01010000;
#1 $display("%b", po);
#1 pi=8'b01010001;
#1 $display("%b", po);
#1 pi=8'b01010010;
#1 $display("%b", po);
#1 pi=8'b01010011;
#1 $display("%b", po);
#1 pi=8'b01010100;
#1 $display("%b", po);
#1 pi=8'b01010101;
#1 $display("%b", po);
#1 pi=8'b01010110;
#1 $display("%b", po);
#1 pi=8'b01010111;
#1 $display("%b", po);
#1 pi=8'b01011000;
#1 $display("%b", po);
#1 pi=8'b01011001;
#1 $display("%b", po);
#1 pi=8'b01011010;
#1 $display("%b", po);
#1 pi=8'b01011011;
#1 $display("%b", po);
#1 pi=8'b01011100;
#1 $display("%b", po);
#1 pi=8'b01011101;
#1 $display("%b", po);
#1 pi=8'b01011110;
#1 $display("%b", po);
#1 pi=8'b01011111;
#1 $display("%b", po);
#1 pi=8'b01100000;
#1 $display("%b", po);
#1 pi=8'b01100001;
#1 $display("%b", po);
#1 pi=8'b01100010;
#1 $display("%b", po);
#1 pi=8'b01100011;
#1 $display("%b", po);
end
endmodule
